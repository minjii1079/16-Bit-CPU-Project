LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY modified_dec3to8 IS
    PORT (
        w  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        En : IN  STD_LOGIC;                   
        y  : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END modified_dec3to8;

ARCHITECTURE Behavior OF modified_dec3to8 IS
    SIGNAL Enw: STD_LOGIC_VECTOR(4 DOWNTO 0); 
BEGIN
    Enw <= En & w;

    WITH Enw SELECT							-- Functions
		y <= 	"0000000000000001" WHEN "10000", --1
				"0000000000000010" WHEN "10001", --2
				"0000000000000100" WHEN "10010", --3
				"0000000000001000" WHEN "10011", --4
				"0000000000010000" WHEN "10100", --5
				"0000000000100000" WHEN "10101", --6
				"0000000001000000" WHEN "10110", --7
				"0000000010000000" WHEN "10111", --8
				"0000000000000000" WHEN OTHERS;
END Behavior;
