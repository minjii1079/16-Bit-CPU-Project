LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;

entity ALU_unit2 is -- ALU unit includes Reg. 3
port ( clk : in std_logic ;
opcode : in std_logic_vector(15 downto 0); -- 8-bit opcode from Decoder
  A, B : inout std_logic_vector(7 downto 0);
neg : out std_logic;
R1, R2 : out std_logic_vector(3 downto 0));  -- R1 = A, R2 = B
end ALU_unit2 ;

architecture calculation of ALU_unit2 is
SIGNAL Result, Reg1, Reg2: std_logic_vector(7 downto 0); -- 8-bit Result
--Reg1, Reg2, 

begin
--Reg1 <= A;
--Reg2 <= B;
process (clk)
begin
if (clk'EVENT AND clk = '1') then
neg <= '0';
case opcode is
when "0000000000000001" => 
     Result(7) <= A(0);
     Result(6) <= A(1);
     Result(5) <= A(2);
     Result(4) <= A(3);
     Result(3) <= A(4);
     Result(2) <= A(5);
     Result(1) <= A(6);
     Result(0) <= A(7);
when "0000000000000010" => 
	Result(7) <= A(7);
	Result(6) <= A(6);
	Result(5) <= A(5);
	Result(4) <= A(4);
	Result(3 downto 0) <= "1111";
when "0000000000000100" =>
Result <= B;
Result(7) <= NOT B(7);
Result(6) <= NOT B(6);
Result(5) <= NOT B(5);
Result(4) <= NOT B(4);
when "0000000000001000" => 
if (A < B) then
Result <= A;
else
Result <= B;
end if;
when "0000000000010000" => 
Result <= (A + B) + 4;
when "0000000000100000" => 
Result <= A + 3;
when "0000000001000000" => 
Result <= A;
Result(0) <= B(0);  --Replace the even bits of A with even bits of B
Result(2) <= B(2);
Result(4) <= B(4);
Result(6) <= B(6);
when "0000000010000000" => 
Result <= NOT(A XOR B);  -- XNORing A and B
when others =>
-- Dont care, do nothing
end case;
end if;
end process;
R1 <= Result(7 DOWNTO 4);
R2 <= Result(3 DOWNTO 0);
end calculation;